`define CLOCK_PERIOD 1.0
