VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SRAM1RW32x50
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN SRAM1RW32x50 0 0 ;
  SIZE 112.368 BY 104.064 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.528 112.368 6.912 ;
        RECT 0.0 14.208 112.368 14.592 ;
        RECT 0.0 21.888 112.368 22.272 ;
        RECT 0.0 29.568 112.368 29.952 ;
        RECT 0.0 37.248 112.368 37.632 ;
        RECT 0.0 44.928 112.368 45.312 ;
        RECT 0.0 52.608 112.368 52.992 ;
        RECT 0.0 60.288 112.368 60.672 ;
        RECT 0.0 67.968 112.368 68.352 ;
        RECT 0.0 75.648 112.368 76.032 ;
        RECT 0.0 83.328 112.368 83.712 ;
        RECT 0.0 91.008 112.368 91.392 ;
        RECT 0.0 98.688 112.368 99.072 ;
    END 
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.296 112.368 7.68 ;
        RECT 0.0 14.976 112.368 15.36 ;
        RECT 0.0 22.656 112.368 23.04 ;
        RECT 0.0 30.336 112.368 30.72 ;
        RECT 0.0 38.016 112.368 38.4 ;
        RECT 0.0 45.696 112.368 46.08 ;
        RECT 0.0 53.376 112.368 53.76 ;
        RECT 0.0 61.056 112.368 61.44 ;
        RECT 0.0 68.736 112.368 69.12 ;
        RECT 0.0 76.416 112.368 76.8 ;
        RECT 0.0 84.096 112.368 84.48 ;
        RECT 0.0 91.776 112.368 92.16 ;
        RECT 0.0 99.456 112.368 99.84 ;
    END 
  END VSS
  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.536 16.0 3.072 ;
    END 
  END CE
  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.608 16.0 6.144 ;
    END 
  END WEB
  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.68 16.0 9.216 ;
    END 
  END OEB
  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.752 16.0 12.288 ;
    END 
  END CSB
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.824 16.0 15.36 ;
    END 
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.896 16.0 18.432 ;
    END 
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.968 16.0 21.504 ;
    END 
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.04 16.0 24.576 ;
    END 
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 32.256 16.0 33.792 ;
    END 
  END A[4]
  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 35.328 16.0 36.864 ;
    END 
  END I[0]
  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 38.4 16.0 39.936 ;
    END 
  END I[1]
  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 41.472 16.0 43.008 ;
    END 
  END I[2]
  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 44.544 16.0 46.08 ;
    END 
  END I[3]
  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 47.616 16.0 49.152 ;
    END 
  END I[4]
  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 50.688 16.0 52.224 ;
    END 
  END I[5]
  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 53.76 16.0 55.296 ;
    END 
  END I[6]
  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 62.976 16.0 64.512 ;
    END 
  END I[7]
  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 66.048 16.0 67.584 ;
    END 
  END I[8]
  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 69.12 16.0 70.656 ;
    END 
  END I[9]
  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 72.192 16.0 73.728 ;
    END 
  END I[10]
  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 75.264 16.0 76.8 ;
    END 
  END I[11]
  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 78.336 16.0 79.872 ;
    END 
  END I[12]
  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 81.408 16.0 82.944 ;
    END 
  END I[13]
  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 84.48 16.0 86.016 ;
    END 
  END I[14]
  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 93.696 16.0 95.232 ;
    END 
  END I[15]
  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 96.768 16.0 98.304 ;
    END 
  END I[16]
  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 99.84 16.0 101.376 ;
    END 
  END I[17]
  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 102.912 16.0 104.448 ;
    END 
  END I[18]
  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 105.984 16.0 107.52 ;
    END 
  END I[19]
  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 109.056 16.0 110.592 ;
    END 
  END I[20]
  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 112.128 16.0 113.664 ;
    END 
  END I[21]
  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 115.2 16.0 116.736 ;
    END 
  END I[22]
  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 124.416 16.0 125.952 ;
    END 
  END I[23]
  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 127.488 16.0 129.024 ;
    END 
  END I[24]
  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 130.56 16.0 132.096 ;
    END 
  END I[25]
  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 133.632 16.0 135.168 ;
    END 
  END I[26]
  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 136.704 16.0 138.24 ;
    END 
  END I[27]
  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 139.776 16.0 141.312 ;
    END 
  END I[28]
  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 142.848 16.0 144.384 ;
    END 
  END I[29]
  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 145.92 16.0 147.456 ;
    END 
  END I[30]
  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 155.136 16.0 156.672 ;
    END 
  END I[31]
  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 158.208 16.0 159.744 ;
    END 
  END I[32]
  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 161.28 16.0 162.816 ;
    END 
  END I[33]
  PIN I[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 164.352 16.0 165.888 ;
    END 
  END I[34]
  PIN I[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 167.424 16.0 168.96 ;
    END 
  END I[35]
  PIN I[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 170.496 16.0 172.032 ;
    END 
  END I[36]
  PIN I[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 173.568 16.0 175.104 ;
    END 
  END I[37]
  PIN I[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 176.64 16.0 178.176 ;
    END 
  END I[38]
  PIN I[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 185.856 16.0 187.392 ;
    END 
  END I[39]
  PIN I[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 188.928 16.0 190.464 ;
    END 
  END I[40]
  PIN I[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 192.0 16.0 193.536 ;
    END 
  END I[41]
  PIN I[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 195.072 16.0 196.608 ;
    END 
  END I[42]
  PIN I[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 198.144 16.0 199.68 ;
    END 
  END I[43]
  PIN I[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 201.216 16.0 202.752 ;
    END 
  END I[44]
  PIN I[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 204.288 16.0 205.824 ;
    END 
  END I[45]
  PIN I[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 207.36 16.0 208.896 ;
    END 
  END I[46]
  PIN I[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 216.576 16.0 218.112 ;
    END 
  END I[47]
  PIN I[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 219.648 16.0 221.184 ;
    END 
  END I[48]
  PIN I[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 222.72 16.0 224.256 ;
    END 
  END I[49]
  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 225.792 16.0 227.328 ;
    END 
  END O[0]
  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 228.864 16.0 230.4 ;
    END 
  END O[1]
  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 231.936 16.0 233.472 ;
    END 
  END O[2]
  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 235.008 16.0 236.544 ;
    END 
  END O[3]
  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 238.08 16.0 239.616 ;
    END 
  END O[4]
  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 247.296 16.0 248.832 ;
    END 
  END O[5]
  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 250.368 16.0 251.904 ;
    END 
  END O[6]
  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 253.44 16.0 254.976 ;
    END 
  END O[7]
  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 256.512 16.0 258.048 ;
    END 
  END O[8]
  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 259.584 16.0 261.12 ;
    END 
  END O[9]
  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 262.656 16.0 264.192 ;
    END 
  END O[10]
  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 265.728 16.0 267.264 ;
    END 
  END O[11]
  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 268.8 16.0 270.336 ;
    END 
  END O[12]
  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 278.016 16.0 279.552 ;
    END 
  END O[13]
  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 281.088 16.0 282.624 ;
    END 
  END O[14]
  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 284.16 16.0 285.696 ;
    END 
  END O[15]
  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 287.232 16.0 288.768 ;
    END 
  END O[16]
  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 290.304 16.0 291.84 ;
    END 
  END O[17]
  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 293.376 16.0 294.912 ;
    END 
  END O[18]
  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 296.448 16.0 297.984 ;
    END 
  END O[19]
  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 299.52 16.0 301.056 ;
    END 
  END O[20]
  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 308.736 16.0 310.272 ;
    END 
  END O[21]
  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 311.808 16.0 313.344 ;
    END 
  END O[22]
  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 314.88 16.0 316.416 ;
    END 
  END O[23]
  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 317.952 16.0 319.488 ;
    END 
  END O[24]
  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 321.024 16.0 322.56 ;
    END 
  END O[25]
  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 324.096 16.0 325.632 ;
    END 
  END O[26]
  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 327.168 16.0 328.704 ;
    END 
  END O[27]
  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 330.24 16.0 331.776 ;
    END 
  END O[28]
  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 333.312 16.0 334.848 ;
    END 
  END O[29]
  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 339.456 16.0 340.992 ;
    END 
  END O[30]
  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 342.528 16.0 344.064 ;
    END 
  END O[31]
  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 345.6 16.0 347.136 ;
    END 
  END O[32]
  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 348.672 16.0 350.208 ;
    END 
  END O[33]
  PIN O[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 351.744 16.0 353.28 ;
    END 
  END O[34]
  PIN O[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 354.816 16.0 356.352 ;
    END 
  END O[35]
  PIN O[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 357.888 16.0 359.424 ;
    END 
  END O[36]
  PIN O[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 360.96 16.0 362.496 ;
    END 
  END O[37]
  PIN O[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 370.176 16.0 371.712 ;
    END 
  END O[38]
  PIN O[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 373.248 16.0 374.784 ;
    END 
  END O[39]
  PIN O[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 376.32 16.0 377.856 ;
    END 
  END O[40]
  PIN O[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 379.392 16.0 380.928 ;
    END 
  END O[41]
  PIN O[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 382.464 16.0 384.0 ;
    END 
  END O[42]
  PIN O[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 385.536 16.0 387.072 ;
    END 
  END O[43]
  PIN O[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 388.608 16.0 390.144 ;
    END 
  END O[44]
  PIN O[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 391.68 16.0 393.216 ;
    END 
  END O[45]
  PIN O[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 400.896 16.0 402.432 ;
    END 
  END O[46]
  PIN O[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 403.968 16.0 405.504 ;
    END 
  END O[47]
  PIN O[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 407.04 16.0 408.576 ;
    END 
  END O[48]
  PIN O[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 410.112 16.0 411.648 ;
    END 
  END O[49]
  OBS 
    LAYER M1 ;
      RECT 4.0 0.0 112.368 104.064 ;
    LAYER M2 ;
      RECT 4.0 0.0 112.368 104.064 ;
    LAYER M3 ;
      RECT 4.0 0.0 112.368 104.064 ;
  END 
END SRAM1RW32x50

END LIBRARY