VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SRAM2RW64x32
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN SRAM2RW64x32 0 0 ;
  SIZE 20.0 BY 141.696 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.528 20.0 6.912 ;
        RECT 0.0 14.208 20.0 14.592 ;
        RECT 0.0 21.888 20.0 22.272 ;
        RECT 0.0 29.568 20.0 29.952 ;
        RECT 0.0 37.248 20.0 37.632 ;
        RECT 0.0 44.928 20.0 45.312 ;
        RECT 0.0 52.608 20.0 52.992 ;
        RECT 0.0 60.288 20.0 60.672 ;
        RECT 0.0 67.968 20.0 68.352 ;
        RECT 0.0 75.648 20.0 76.032 ;
        RECT 0.0 83.328 20.0 83.712 ;
        RECT 0.0 91.008 20.0 91.392 ;
        RECT 0.0 98.688 20.0 99.072 ;
        RECT 0.0 106.368 20.0 106.752 ;
        RECT 0.0 114.048 20.0 114.432 ;
        RECT 0.0 121.728 20.0 122.112 ;
        RECT 0.0 129.408 20.0 129.792 ;
        RECT 0.0 137.088 20.0 137.472 ;
    END 
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.296 20.0 7.68 ;
        RECT 0.0 14.976 20.0 15.36 ;
        RECT 0.0 22.656 20.0 23.04 ;
        RECT 0.0 30.336 20.0 30.72 ;
        RECT 0.0 38.016 20.0 38.4 ;
        RECT 0.0 45.696 20.0 46.08 ;
        RECT 0.0 53.376 20.0 53.76 ;
        RECT 0.0 61.056 20.0 61.44 ;
        RECT 0.0 68.736 20.0 69.12 ;
        RECT 0.0 76.416 20.0 76.8 ;
        RECT 0.0 84.096 20.0 84.48 ;
        RECT 0.0 91.776 20.0 92.16 ;
        RECT 0.0 99.456 20.0 99.84 ;
        RECT 0.0 107.136 20.0 107.52 ;
        RECT 0.0 114.816 20.0 115.2 ;
        RECT 0.0 122.496 20.0 122.88 ;
        RECT 0.0 130.176 20.0 130.56 ;
        RECT 0.0 137.856 20.0 138.24 ;
    END 
  END VSS
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.384 4.0 0.768 ;
    END 
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.152 4.0 1.536 ;
    END 
  END CE2
  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.92 4.0 2.304 ;
    END 
  END WEB1
  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.688 4.0 3.072 ;
    END 
  END WEB2
  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 3.456 4.0 3.84 ;
    END 
  END OEB1
  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.224 4.0 4.608 ;
    END 
  END OEB2
  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.992 4.0 5.376 ;
    END 
  END CSB1
  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 5.76 4.0 6.144 ;
    END 
  END CSB2
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.064 4.0 8.448 ;
    END 
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.832 4.0 9.216 ;
    END 
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 9.6 4.0 9.984 ;
    END 
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.368 4.0 10.752 ;
    END 
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.136 4.0 11.52 ;
    END 
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.904 4.0 12.288 ;
    END 
  END A1[5]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.672 4.0 13.056 ;
    END 
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.44 4.0 13.824 ;
    END 
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 15.744 4.0 16.128 ;
    END 
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.512 4.0 16.896 ;
    END 
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.28 4.0 17.664 ;
    END 
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.048 4.0 18.432 ;
    END 
  END A2[5]
  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.816 4.0 19.2 ;
    END 
  END I1[0]
  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.584 4.0 19.968 ;
    END 
  END I1[1]
  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 20.352 4.0 20.736 ;
    END 
  END I1[2]
  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.12 4.0 21.504 ;
    END 
  END I1[3]
  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.424 4.0 23.808 ;
    END 
  END I1[4]
  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.192 4.0 24.576 ;
    END 
  END I1[5]
  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.96 4.0 25.344 ;
    END 
  END I1[6]
  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.728 4.0 26.112 ;
    END 
  END I1[7]
  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 26.496 4.0 26.88 ;
    END 
  END I1[8]
  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 27.264 4.0 27.648 ;
    END 
  END I1[9]
  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 28.032 4.0 28.416 ;
    END 
  END I1[10]
  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 28.8 4.0 29.184 ;
    END 
  END I1[11]
  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.104 4.0 31.488 ;
    END 
  END I1[12]
  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.872 4.0 32.256 ;
    END 
  END I1[13]
  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 32.64 4.0 33.024 ;
    END 
  END I1[14]
  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 33.408 4.0 33.792 ;
    END 
  END I1[15]
  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 34.176 4.0 34.56 ;
    END 
  END I1[16]
  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 34.944 4.0 35.328 ;
    END 
  END I1[17]
  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 35.712 4.0 36.096 ;
    END 
  END I1[18]
  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 36.48 4.0 36.864 ;
    END 
  END I1[19]
  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 38.784 4.0 39.168 ;
    END 
  END I1[20]
  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 39.552 4.0 39.936 ;
    END 
  END I1[21]
  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 40.32 4.0 40.704 ;
    END 
  END I1[22]
  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 41.088 4.0 41.472 ;
    END 
  END I1[23]
  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 41.856 4.0 42.24 ;
    END 
  END I1[24]
  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 42.624 4.0 43.008 ;
    END 
  END I1[25]
  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 43.392 4.0 43.776 ;
    END 
  END I1[26]
  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 44.16 4.0 44.544 ;
    END 
  END I1[27]
  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 46.464 4.0 46.848 ;
    END 
  END I1[28]
  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 47.232 4.0 47.616 ;
    END 
  END I1[29]
  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 48.0 4.0 48.384 ;
    END 
  END I1[30]
  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 48.768 4.0 49.152 ;
    END 
  END I1[31]
  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 49.536 4.0 49.92 ;
    END 
  END I2[0]
  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 50.304 4.0 50.688 ;
    END 
  END I2[1]
  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 51.072 4.0 51.456 ;
    END 
  END I2[2]
  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 51.84 4.0 52.224 ;
    END 
  END I2[3]
  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 54.144 4.0 54.528 ;
    END 
  END I2[4]
  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 54.912 4.0 55.296 ;
    END 
  END I2[5]
  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 55.68 4.0 56.064 ;
    END 
  END I2[6]
  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 56.448 4.0 56.832 ;
    END 
  END I2[7]
  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 57.216 4.0 57.6 ;
    END 
  END I2[8]
  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 57.984 4.0 58.368 ;
    END 
  END I2[9]
  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 58.752 4.0 59.136 ;
    END 
  END I2[10]
  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 59.52 4.0 59.904 ;
    END 
  END I2[11]
  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 61.824 4.0 62.208 ;
    END 
  END I2[12]
  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 62.592 4.0 62.976 ;
    END 
  END I2[13]
  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 63.36 4.0 63.744 ;
    END 
  END I2[14]
  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 64.128 4.0 64.512 ;
    END 
  END I2[15]
  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 64.896 4.0 65.28 ;
    END 
  END I2[16]
  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 65.664 4.0 66.048 ;
    END 
  END I2[17]
  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 66.432 4.0 66.816 ;
    END 
  END I2[18]
  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 67.2 4.0 67.584 ;
    END 
  END I2[19]
  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 69.504 4.0 69.888 ;
    END 
  END I2[20]
  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 70.272 4.0 70.656 ;
    END 
  END I2[21]
  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 71.04 4.0 71.424 ;
    END 
  END I2[22]
  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 71.808 4.0 72.192 ;
    END 
  END I2[23]
  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 72.576 4.0 72.96 ;
    END 
  END I2[24]
  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 73.344 4.0 73.728 ;
    END 
  END I2[25]
  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 74.112 4.0 74.496 ;
    END 
  END I2[26]
  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 74.88 4.0 75.264 ;
    END 
  END I2[27]
  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 77.184 4.0 77.568 ;
    END 
  END I2[28]
  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 77.952 4.0 78.336 ;
    END 
  END I2[29]
  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 78.72 4.0 79.104 ;
    END 
  END I2[30]
  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 79.488 4.0 79.872 ;
    END 
  END I2[31]
  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 80.256 4.0 80.64 ;
    END 
  END O1[0]
  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 81.024 4.0 81.408 ;
    END 
  END O1[1]
  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 81.792 4.0 82.176 ;
    END 
  END O1[2]
  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 82.56 4.0 82.944 ;
    END 
  END O1[3]
  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 84.864 4.0 85.248 ;
    END 
  END O1[4]
  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 85.632 4.0 86.016 ;
    END 
  END O1[5]
  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 86.4 4.0 86.784 ;
    END 
  END O1[6]
  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 87.168 4.0 87.552 ;
    END 
  END O1[7]
  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 87.936 4.0 88.32 ;
    END 
  END O1[8]
  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 88.704 4.0 89.088 ;
    END 
  END O1[9]
  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 89.472 4.0 89.856 ;
    END 
  END O1[10]
  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 90.24 4.0 90.624 ;
    END 
  END O1[11]
  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 92.544 4.0 92.928 ;
    END 
  END O1[12]
  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 93.312 4.0 93.696 ;
    END 
  END O1[13]
  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 94.08 4.0 94.464 ;
    END 
  END O1[14]
  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 94.848 4.0 95.232 ;
    END 
  END O1[15]
  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 95.616 4.0 96.0 ;
    END 
  END O1[16]
  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 96.384 4.0 96.768 ;
    END 
  END O1[17]
  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 97.152 4.0 97.536 ;
    END 
  END O1[18]
  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 97.92 4.0 98.304 ;
    END 
  END O1[19]
  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 100.224 4.0 100.608 ;
    END 
  END O1[20]
  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 100.992 4.0 101.376 ;
    END 
  END O1[21]
  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 101.76 4.0 102.144 ;
    END 
  END O1[22]
  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 102.528 4.0 102.912 ;
    END 
  END O1[23]
  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 103.296 4.0 103.68 ;
    END 
  END O1[24]
  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 104.064 4.0 104.448 ;
    END 
  END O1[25]
  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 104.832 4.0 105.216 ;
    END 
  END O1[26]
  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 105.6 4.0 105.984 ;
    END 
  END O1[27]
  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 107.904 4.0 108.288 ;
    END 
  END O1[28]
  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 108.672 4.0 109.056 ;
    END 
  END O1[29]
  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 109.44 4.0 109.824 ;
    END 
  END O1[30]
  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 110.208 4.0 110.592 ;
    END 
  END O1[31]
  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 110.976 4.0 111.36 ;
    END 
  END O2[0]
  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 111.744 4.0 112.128 ;
    END 
  END O2[1]
  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 112.512 4.0 112.896 ;
    END 
  END O2[2]
  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 113.28 4.0 113.664 ;
    END 
  END O2[3]
  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 115.584 4.0 115.968 ;
    END 
  END O2[4]
  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 116.352 4.0 116.736 ;
    END 
  END O2[5]
  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 117.12 4.0 117.504 ;
    END 
  END O2[6]
  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 117.888 4.0 118.272 ;
    END 
  END O2[7]
  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 118.656 4.0 119.04 ;
    END 
  END O2[8]
  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 119.424 4.0 119.808 ;
    END 
  END O2[9]
  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 120.192 4.0 120.576 ;
    END 
  END O2[10]
  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 120.96 4.0 121.344 ;
    END 
  END O2[11]
  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 123.264 4.0 123.648 ;
    END 
  END O2[12]
  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 124.032 4.0 124.416 ;
    END 
  END O2[13]
  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 124.8 4.0 125.184 ;
    END 
  END O2[14]
  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 125.568 4.0 125.952 ;
    END 
  END O2[15]
  PIN O2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 126.336 4.0 126.72 ;
    END 
  END O2[16]
  PIN O2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 127.104 4.0 127.488 ;
    END 
  END O2[17]
  PIN O2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 127.872 4.0 128.256 ;
    END 
  END O2[18]
  PIN O2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 128.64 4.0 129.024 ;
    END 
  END O2[19]
  PIN O2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 130.944 4.0 131.328 ;
    END 
  END O2[20]
  PIN O2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 131.712 4.0 132.096 ;
    END 
  END O2[21]
  PIN O2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 132.48 4.0 132.864 ;
    END 
  END O2[22]
  PIN O2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 133.248 4.0 133.632 ;
    END 
  END O2[23]
  PIN O2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 134.016 4.0 134.4 ;
    END 
  END O2[24]
  PIN O2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 134.784 4.0 135.168 ;
    END 
  END O2[25]
  PIN O2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 135.552 4.0 135.936 ;
    END 
  END O2[26]
  PIN O2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 136.32 4.0 136.704 ;
    END 
  END O2[27]
  PIN O2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 138.624 4.0 139.008 ;
    END 
  END O2[28]
  PIN O2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 139.392 4.0 139.776 ;
    END 
  END O2[29]
  PIN O2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 140.16 4.0 140.544 ;
    END 
  END O2[30]
  PIN O2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 140.928 4.0 141.312 ;
    END 
  END O2[31]
  OBS 
    LAYER M1 ;
      RECT 4.0 0.0 20.0 141.696 ;
    LAYER M2 ;
      RECT 4.0 0.0 20.0 141.696 ;
    LAYER M3 ;
      RECT 4.0 0.0 20.0 141.696 ;
  END 
END SRAM2RW64x32

END LIBRARY