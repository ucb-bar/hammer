VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SRAM2RW32x33
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN SRAM2RW32x33 0 0 ;
  SIZE 32.928 BY 35.808 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.632 32.928 1.728 ;
        RECT 0.0 3.552 32.928 3.648 ;
        RECT 0.0 5.472 32.928 5.568 ;
        RECT 0.0 7.392 32.928 7.488 ;
        RECT 0.0 9.312 32.928 9.408 ;
        RECT 0.0 11.232 32.928 11.328 ;
        RECT 0.0 13.152 32.928 13.248 ;
        RECT 0.0 15.072 32.928 15.168 ;
        RECT 0.0 16.992 32.928 17.088 ;
        RECT 0.0 18.912 32.928 19.008 ;
        RECT 0.0 20.832 32.928 20.928 ;
        RECT 0.0 22.752 32.928 22.848 ;
        RECT 0.0 24.672 32.928 24.768 ;
        RECT 0.0 26.592 32.928 26.688 ;
        RECT 0.0 28.512 32.928 28.608 ;
        RECT 0.0 30.432 32.928 30.528 ;
        RECT 0.0 32.352 32.928 32.448 ;
        RECT 0.0 34.272 32.928 34.368 ;
    END 
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.824 32.928 1.92 ;
        RECT 0.0 3.744 32.928 3.84 ;
        RECT 0.0 5.664 32.928 5.76 ;
        RECT 0.0 7.584 32.928 7.68 ;
        RECT 0.0 9.504 32.928 9.6 ;
        RECT 0.0 11.424 32.928 11.52 ;
        RECT 0.0 13.344 32.928 13.44 ;
        RECT 0.0 15.264 32.928 15.36 ;
        RECT 0.0 17.184 32.928 17.28 ;
        RECT 0.0 19.104 32.928 19.2 ;
        RECT 0.0 21.024 32.928 21.12 ;
        RECT 0.0 22.944 32.928 23.04 ;
        RECT 0.0 24.864 32.928 24.96 ;
        RECT 0.0 26.784 32.928 26.88 ;
        RECT 0.0 28.704 32.928 28.8 ;
        RECT 0.0 30.624 32.928 30.72 ;
        RECT 0.0 32.544 32.928 32.64 ;
        RECT 0.0 34.464 32.928 34.56 ;
    END 
  END VSS
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.096 4.0 0.192 ;
    END 
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.288 4.0 0.384 ;
    END 
  END CE2
  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.48 4.0 0.576 ;
    END 
  END WEB1
  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.672 4.0 0.768 ;
    END 
  END WEB2
  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.864 4.0 0.96 ;
    END 
  END OEB1
  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.056 4.0 1.152 ;
    END 
  END OEB2
  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.248 4.0 1.344 ;
    END 
  END CSB1
  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.44 4.0 1.536 ;
    END 
  END CSB2
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.016 4.0 2.112 ;
    END 
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.208 4.0 2.304 ;
    END 
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.4 4.0 2.496 ;
    END 
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.592 4.0 2.688 ;
    END 
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.784 4.0 2.88 ;
    END 
  END A1[4]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.976 4.0 3.072 ;
    END 
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 3.168 4.0 3.264 ;
    END 
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 3.36 4.0 3.456 ;
    END 
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 3.936 4.0 4.032 ;
    END 
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.128 4.0 4.224 ;
    END 
  END A2[4]
  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.32 4.0 4.416 ;
    END 
  END I1[0]
  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.512 4.0 4.608 ;
    END 
  END I1[1]
  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.704 4.0 4.8 ;
    END 
  END I1[2]
  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.896 4.0 4.992 ;
    END 
  END I1[3]
  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 5.088 4.0 5.184 ;
    END 
  END I1[4]
  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 5.28 4.0 5.376 ;
    END 
  END I1[5]
  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 5.856 4.0 5.952 ;
    END 
  END I1[6]
  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.048 4.0 6.144 ;
    END 
  END I1[7]
  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.24 4.0 6.336 ;
    END 
  END I1[8]
  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.432 4.0 6.528 ;
    END 
  END I1[9]
  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.624 4.0 6.72 ;
    END 
  END I1[10]
  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.816 4.0 6.912 ;
    END 
  END I1[11]
  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.008 4.0 7.104 ;
    END 
  END I1[12]
  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.2 4.0 7.296 ;
    END 
  END I1[13]
  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.776 4.0 7.872 ;
    END 
  END I1[14]
  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.968 4.0 8.064 ;
    END 
  END I1[15]
  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.16 4.0 8.256 ;
    END 
  END I1[16]
  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.352 4.0 8.448 ;
    END 
  END I1[17]
  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.544 4.0 8.64 ;
    END 
  END I1[18]
  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.736 4.0 8.832 ;
    END 
  END I1[19]
  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.928 4.0 9.024 ;
    END 
  END I1[20]
  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 9.12 4.0 9.216 ;
    END 
  END I1[21]
  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 9.696 4.0 9.792 ;
    END 
  END I1[22]
  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 9.888 4.0 9.984 ;
    END 
  END I1[23]
  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.08 4.0 10.176 ;
    END 
  END I1[24]
  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.272 4.0 10.368 ;
    END 
  END I1[25]
  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.464 4.0 10.56 ;
    END 
  END I1[26]
  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.656 4.0 10.752 ;
    END 
  END I1[27]
  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.848 4.0 10.944 ;
    END 
  END I1[28]
  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.04 4.0 11.136 ;
    END 
  END I1[29]
  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.616 4.0 11.712 ;
    END 
  END I1[30]
  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.808 4.0 11.904 ;
    END 
  END I1[31]
  PIN I1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.0 4.0 12.096 ;
    END 
  END I1[32]
  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.192 4.0 12.288 ;
    END 
  END I2[0]
  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.384 4.0 12.48 ;
    END 
  END I2[1]
  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.576 4.0 12.672 ;
    END 
  END I2[2]
  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.768 4.0 12.864 ;
    END 
  END I2[3]
  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.96 4.0 13.056 ;
    END 
  END I2[4]
  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.536 4.0 13.632 ;
    END 
  END I2[5]
  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.728 4.0 13.824 ;
    END 
  END I2[6]
  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.92 4.0 14.016 ;
    END 
  END I2[7]
  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.112 4.0 14.208 ;
    END 
  END I2[8]
  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.304 4.0 14.4 ;
    END 
  END I2[9]
  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.496 4.0 14.592 ;
    END 
  END I2[10]
  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.688 4.0 14.784 ;
    END 
  END I2[11]
  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.88 4.0 14.976 ;
    END 
  END I2[12]
  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 15.456 4.0 15.552 ;
    END 
  END I2[13]
  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 15.648 4.0 15.744 ;
    END 
  END I2[14]
  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 15.84 4.0 15.936 ;
    END 
  END I2[15]
  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.032 4.0 16.128 ;
    END 
  END I2[16]
  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.224 4.0 16.32 ;
    END 
  END I2[17]
  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.416 4.0 16.512 ;
    END 
  END I2[18]
  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.608 4.0 16.704 ;
    END 
  END I2[19]
  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.8 4.0 16.896 ;
    END 
  END I2[20]
  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.376 4.0 17.472 ;
    END 
  END I2[21]
  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.568 4.0 17.664 ;
    END 
  END I2[22]
  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.76 4.0 17.856 ;
    END 
  END I2[23]
  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.952 4.0 18.048 ;
    END 
  END I2[24]
  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.144 4.0 18.24 ;
    END 
  END I2[25]
  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.336 4.0 18.432 ;
    END 
  END I2[26]
  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.528 4.0 18.624 ;
    END 
  END I2[27]
  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.72 4.0 18.816 ;
    END 
  END I2[28]
  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.296 4.0 19.392 ;
    END 
  END I2[29]
  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.488 4.0 19.584 ;
    END 
  END I2[30]
  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.68 4.0 19.776 ;
    END 
  END I2[31]
  PIN I2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.872 4.0 19.968 ;
    END 
  END I2[32]
  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 20.064 4.0 20.16 ;
    END 
  END O1[0]
  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 20.256 4.0 20.352 ;
    END 
  END O1[1]
  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 20.448 4.0 20.544 ;
    END 
  END O1[2]
  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 20.64 4.0 20.736 ;
    END 
  END O1[3]
  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.216 4.0 21.312 ;
    END 
  END O1[4]
  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.408 4.0 21.504 ;
    END 
  END O1[5]
  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.6 4.0 21.696 ;
    END 
  END O1[6]
  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.792 4.0 21.888 ;
    END 
  END O1[7]
  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.984 4.0 22.08 ;
    END 
  END O1[8]
  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 22.176 4.0 22.272 ;
    END 
  END O1[9]
  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 22.368 4.0 22.464 ;
    END 
  END O1[10]
  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 22.56 4.0 22.656 ;
    END 
  END O1[11]
  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.136 4.0 23.232 ;
    END 
  END O1[12]
  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.328 4.0 23.424 ;
    END 
  END O1[13]
  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.52 4.0 23.616 ;
    END 
  END O1[14]
  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.712 4.0 23.808 ;
    END 
  END O1[15]
  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.904 4.0 24.0 ;
    END 
  END O1[16]
  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.096 4.0 24.192 ;
    END 
  END O1[17]
  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.288 4.0 24.384 ;
    END 
  END O1[18]
  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.48 4.0 24.576 ;
    END 
  END O1[19]
  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.056 4.0 25.152 ;
    END 
  END O1[20]
  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.248 4.0 25.344 ;
    END 
  END O1[21]
  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.44 4.0 25.536 ;
    END 
  END O1[22]
  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.632 4.0 25.728 ;
    END 
  END O1[23]
  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.824 4.0 25.92 ;
    END 
  END O1[24]
  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 26.016 4.0 26.112 ;
    END 
  END O1[25]
  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 26.208 4.0 26.304 ;
    END 
  END O1[26]
  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 26.4 4.0 26.496 ;
    END 
  END O1[27]
  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 26.976 4.0 27.072 ;
    END 
  END O1[28]
  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 27.168 4.0 27.264 ;
    END 
  END O1[29]
  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 27.36 4.0 27.456 ;
    END 
  END O1[30]
  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 27.552 4.0 27.648 ;
    END 
  END O1[31]
  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 27.744 4.0 27.84 ;
    END 
  END O1[32]
  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 27.936 4.0 28.032 ;
    END 
  END O2[0]
  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 28.128 4.0 28.224 ;
    END 
  END O2[1]
  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 28.32 4.0 28.416 ;
    END 
  END O2[2]
  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 28.896 4.0 28.992 ;
    END 
  END O2[3]
  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 29.088 4.0 29.184 ;
    END 
  END O2[4]
  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 29.28 4.0 29.376 ;
    END 
  END O2[5]
  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 29.472 4.0 29.568 ;
    END 
  END O2[6]
  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 29.664 4.0 29.76 ;
    END 
  END O2[7]
  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 29.856 4.0 29.952 ;
    END 
  END O2[8]
  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 30.048 4.0 30.144 ;
    END 
  END O2[9]
  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 30.24 4.0 30.336 ;
    END 
  END O2[10]
  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 30.816 4.0 30.912 ;
    END 
  END O2[11]
  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.008 4.0 31.104 ;
    END 
  END O2[12]
  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.2 4.0 31.296 ;
    END 
  END O2[13]
  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.392 4.0 31.488 ;
    END 
  END O2[14]
  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.584 4.0 31.68 ;
    END 
  END O2[15]
  PIN O2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.776 4.0 31.872 ;
    END 
  END O2[16]
  PIN O2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 31.968 4.0 32.064 ;
    END 
  END O2[17]
  PIN O2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 32.16 4.0 32.256 ;
    END 
  END O2[18]
  PIN O2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 32.736 4.0 32.832 ;
    END 
  END O2[19]
  PIN O2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 32.928 4.0 33.024 ;
    END 
  END O2[20]
  PIN O2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 33.12 4.0 33.216 ;
    END 
  END O2[21]
  PIN O2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 33.312 4.0 33.408 ;
    END 
  END O2[22]
  PIN O2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 33.504 4.0 33.6 ;
    END 
  END O2[23]
  PIN O2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 33.696 4.0 33.792 ;
    END 
  END O2[24]
  PIN O2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 33.888 4.0 33.984 ;
    END 
  END O2[25]
  PIN O2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 34.08 4.0 34.176 ;
    END 
  END O2[26]
  PIN O2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 34.656 4.0 34.752 ;
    END 
  END O2[27]
  PIN O2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 34.848 4.0 34.944 ;
    END 
  END O2[28]
  PIN O2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 35.04 4.0 35.136 ;
    END 
  END O2[29]
  PIN O2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 35.232 4.0 35.328 ;
    END 
  END O2[30]
  PIN O2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 35.424 4.0 35.52 ;
    END 
  END O2[31]
  PIN O2[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 35.616 4.0 35.712 ;
    END 
  END O2[32]
  OBS 
    LAYER M1 ;
      RECT 4.0 0.0 32.928 35.808 ;
    LAYER M2 ;
      RECT 4.0 0.0 32.928 35.808 ;
    LAYER M3 ;
      RECT 4.0 0.0 32.928 35.808 ;
  END 
END SRAM2RW32x33

END LIBRARY