`define CLOCK_PERIOD 1.0
`define PRINTF_COND TestDriver.printf_cond
`define STOP_COND !TestDriver.reset
`define RANDOMIZE_MEM_INIT
`define RANDOMIZE_REG_INIT
`define RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE_INVALID_ASSIGN
