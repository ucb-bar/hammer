VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SRAM2RW32x22
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN SRAM2RW32x22 0 0 ;
  SIZE 24.128 BY 28.264 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.632 24.128 1.728 ;
        RECT 0.0 3.552 24.128 3.648 ;
        RECT 0.0 5.472 24.128 5.568 ;
        RECT 0.0 7.392 24.128 7.488 ;
        RECT 0.0 9.312 24.128 9.408 ;
        RECT 0.0 11.232 24.128 11.328 ;
        RECT 0.0 13.152 24.128 13.248 ;
        RECT 0.0 15.072 24.128 15.168 ;
        RECT 0.0 16.992 24.128 17.088 ;
        RECT 0.0 18.912 24.128 19.008 ;
        RECT 0.0 20.832 24.128 20.928 ;
        RECT 0.0 22.752 24.128 22.848 ;
        RECT 0.0 24.672 24.128 24.768 ;
    END 
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.824 24.128 1.92 ;
        RECT 0.0 3.744 24.128 3.84 ;
        RECT 0.0 5.664 24.128 5.76 ;
        RECT 0.0 7.584 24.128 7.68 ;
        RECT 0.0 9.504 24.128 9.6 ;
        RECT 0.0 11.424 24.128 11.52 ;
        RECT 0.0 13.344 24.128 13.44 ;
        RECT 0.0 15.264 24.128 15.36 ;
        RECT 0.0 17.184 24.128 17.28 ;
        RECT 0.0 19.104 24.128 19.2 ;
        RECT 0.0 21.024 24.128 21.12 ;
        RECT 0.0 22.944 24.128 23.04 ;
        RECT 0.0 24.864 24.128 24.96 ;
    END 
  END VSS
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.096 4.0 0.192 ;
    END 
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.288 4.0 0.384 ;
    END 
  END CE2
  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.48 4.0 0.576 ;
    END 
  END WEB1
  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.672 4.0 0.768 ;
    END 
  END WEB2
  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 0.864 4.0 0.96 ;
    END 
  END OEB1
  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.056 4.0 1.152 ;
    END 
  END OEB2
  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.248 4.0 1.344 ;
    END 
  END CSB1
  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 1.44 4.0 1.536 ;
    END 
  END CSB2
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.016 4.0 2.112 ;
    END 
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.208 4.0 2.304 ;
    END 
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.4 4.0 2.496 ;
    END 
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.592 4.0 2.688 ;
    END 
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.784 4.0 2.88 ;
    END 
  END A1[4]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 2.976 4.0 3.072 ;
    END 
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 3.168 4.0 3.264 ;
    END 
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 3.36 4.0 3.456 ;
    END 
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 3.936 4.0 4.032 ;
    END 
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.128 4.0 4.224 ;
    END 
  END A2[4]
  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.32 4.0 4.416 ;
    END 
  END I1[0]
  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.512 4.0 4.608 ;
    END 
  END I1[1]
  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.704 4.0 4.8 ;
    END 
  END I1[2]
  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 4.896 4.0 4.992 ;
    END 
  END I1[3]
  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 5.088 4.0 5.184 ;
    END 
  END I1[4]
  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 5.28 4.0 5.376 ;
    END 
  END I1[5]
  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 5.856 4.0 5.952 ;
    END 
  END I1[6]
  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.048 4.0 6.144 ;
    END 
  END I1[7]
  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.24 4.0 6.336 ;
    END 
  END I1[8]
  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.432 4.0 6.528 ;
    END 
  END I1[9]
  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.624 4.0 6.72 ;
    END 
  END I1[10]
  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 6.816 4.0 6.912 ;
    END 
  END I1[11]
  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.008 4.0 7.104 ;
    END 
  END I1[12]
  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.2 4.0 7.296 ;
    END 
  END I1[13]
  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.776 4.0 7.872 ;
    END 
  END I1[14]
  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 7.968 4.0 8.064 ;
    END 
  END I1[15]
  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.16 4.0 8.256 ;
    END 
  END I1[16]
  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.352 4.0 8.448 ;
    END 
  END I1[17]
  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.544 4.0 8.64 ;
    END 
  END I1[18]
  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.736 4.0 8.832 ;
    END 
  END I1[19]
  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 8.928 4.0 9.024 ;
    END 
  END I1[20]
  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 9.12 4.0 9.216 ;
    END 
  END I1[21]
  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 9.696 4.0 9.792 ;
    END 
  END I2[0]
  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 9.888 4.0 9.984 ;
    END 
  END I2[1]
  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.08 4.0 10.176 ;
    END 
  END I2[2]
  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.272 4.0 10.368 ;
    END 
  END I2[3]
  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.464 4.0 10.56 ;
    END 
  END I2[4]
  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.656 4.0 10.752 ;
    END 
  END I2[5]
  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 10.848 4.0 10.944 ;
    END 
  END I2[6]
  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.04 4.0 11.136 ;
    END 
  END I2[7]
  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.616 4.0 11.712 ;
    END 
  END I2[8]
  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 11.808 4.0 11.904 ;
    END 
  END I2[9]
  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.0 4.0 12.096 ;
    END 
  END I2[10]
  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.192 4.0 12.288 ;
    END 
  END I2[11]
  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.384 4.0 12.48 ;
    END 
  END I2[12]
  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.576 4.0 12.672 ;
    END 
  END I2[13]
  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.768 4.0 12.864 ;
    END 
  END I2[14]
  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 12.96 4.0 13.056 ;
    END 
  END I2[15]
  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.536 4.0 13.632 ;
    END 
  END I2[16]
  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.728 4.0 13.824 ;
    END 
  END I2[17]
  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 13.92 4.0 14.016 ;
    END 
  END I2[18]
  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.112 4.0 14.208 ;
    END 
  END I2[19]
  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.304 4.0 14.4 ;
    END 
  END I2[20]
  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.496 4.0 14.592 ;
    END 
  END I2[21]
  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.688 4.0 14.784 ;
    END 
  END O1[0]
  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 14.88 4.0 14.976 ;
    END 
  END O1[1]
  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 15.456 4.0 15.552 ;
    END 
  END O1[2]
  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 15.648 4.0 15.744 ;
    END 
  END O1[3]
  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 15.84 4.0 15.936 ;
    END 
  END O1[4]
  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.032 4.0 16.128 ;
    END 
  END O1[5]
  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.224 4.0 16.32 ;
    END 
  END O1[6]
  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.416 4.0 16.512 ;
    END 
  END O1[7]
  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.608 4.0 16.704 ;
    END 
  END O1[8]
  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 16.8 4.0 16.896 ;
    END 
  END O1[9]
  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.376 4.0 17.472 ;
    END 
  END O1[10]
  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.568 4.0 17.664 ;
    END 
  END O1[11]
  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.76 4.0 17.856 ;
    END 
  END O1[12]
  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 17.952 4.0 18.048 ;
    END 
  END O1[13]
  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.144 4.0 18.24 ;
    END 
  END O1[14]
  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.336 4.0 18.432 ;
    END 
  END O1[15]
  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.528 4.0 18.624 ;
    END 
  END O1[16]
  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 18.72 4.0 18.816 ;
    END 
  END O1[17]
  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.296 4.0 19.392 ;
    END 
  END O1[18]
  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.488 4.0 19.584 ;
    END 
  END O1[19]
  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.68 4.0 19.776 ;
    END 
  END O1[20]
  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 19.872 4.0 19.968 ;
    END 
  END O1[21]
  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 20.064 4.0 20.16 ;
    END 
  END O2[0]
  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 20.256 4.0 20.352 ;
    END 
  END O2[1]
  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 20.448 4.0 20.544 ;
    END 
  END O2[2]
  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 20.64 4.0 20.736 ;
    END 
  END O2[3]
  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.216 4.0 21.312 ;
    END 
  END O2[4]
  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.408 4.0 21.504 ;
    END 
  END O2[5]
  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.6 4.0 21.696 ;
    END 
  END O2[6]
  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.792 4.0 21.888 ;
    END 
  END O2[7]
  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 21.984 4.0 22.08 ;
    END 
  END O2[8]
  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 22.176 4.0 22.272 ;
    END 
  END O2[9]
  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 22.368 4.0 22.464 ;
    END 
  END O2[10]
  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 22.56 4.0 22.656 ;
    END 
  END O2[11]
  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.136 4.0 23.232 ;
    END 
  END O2[12]
  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.328 4.0 23.424 ;
    END 
  END O2[13]
  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.52 4.0 23.616 ;
    END 
  END O2[14]
  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.712 4.0 23.808 ;
    END 
  END O2[15]
  PIN O2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 23.904 4.0 24.0 ;
    END 
  END O2[16]
  PIN O2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.096 4.0 24.192 ;
    END 
  END O2[17]
  PIN O2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.288 4.0 24.384 ;
    END 
  END O2[18]
  PIN O2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 24.48 4.0 24.576 ;
    END 
  END O2[19]
  PIN O2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.056 4.0 25.152 ;
    END 
  END O2[20]
  PIN O2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.0 25.248 4.0 25.344 ;
    END 
  END O2[21]
  OBS 
    LAYER M1 ;
      RECT 4.0 0.0 24.128 28.264 ;
    LAYER M2 ;
      RECT 4.0 0.0 24.128 28.264 ;
    LAYER M3 ;
      RECT 4.0 0.0 24.128 28.264 ;
  END 
END SRAM2RW32x22

END LIBRARY